`timescale 1ns / 1ps
`include "src/VectorMultiplication.v"

module FloatMultiplicationTB #(parameter VLEN = 5);
    reg [31:0] A, B [0:VLEN-1];  // 5-element float vectors
    wire [(32 * VLEN) - 1:0] A_packed, B_packed;
    reg clk;
    reg overflow, underflow, exception;
    wire [31:0] result;
    real value;  // real (64bit FP) not synthesizable, only for sim comparison

    // pack the A, B arrays
    genvar i;
    for(i = 0; i < VLEN; i = i + 1) begin
        assign A_packed[32 * i +: 31] = A[i];
        assign B_packed[32 * i +: 31] = B[i];
    end

    VectorMultiplication #(.VLEN(VLEN)) mult (.A(A_packed), .B(B_packed), .clk(clk), .result(result));

    // numbers assignments
    initial
    begin
        A[0] = 32'b0_10000000_10011001100110011001100;  // 3.2
        B[0] = 32'b0_10000001_00001100110011001100110;  // 4.2

        A[1] = 32'b0_01111110_01010001111010111000010;  // 0.66
        B[1] = 32'b0_01111110_00000101000111101011100;  // 0.51

        A[2] = 32'b1_01111110_00000000000000000000000;  // -0.5
        B[2] = 32'b1_10000001_10011001100110011001100;  // -6.4

        A[3] = 32'b1_01111110_00000000000000000000000;  // -0.5
        B[3] = 32'b0_10000001_10011001100110011001100;  //  6.4

        A[4] = 32'h4034b4b5;  //  2.82
        B[4] = 32'hbf70f0f1;  // -0.94
    end

    // displaying
    initial
    begin
        // dump to vcd file for GTKWave
        $dumpfile("FloatMultiplicationTb.vcd");
        $dumpvars;

        #100
        value =(2**(result[30:23]-127))*($itor({1'b1,result[22:0]})/2**23)*((-1)**(result[31]));
        $display("Expected Value : %f Result : %f",
                    (3.2 * 4.2) + (0.66 * 0.51) + ((-0.5) * (-6.4)) + ((-0.5) * (6.4)) + (2.82*(-0.94)),
                    value);

        $display("res = %b 1.%b * 2 ^ (%0d - 127)", result[31], result[22:0], result[30:23]);
        $finish;
    end

endmodule
